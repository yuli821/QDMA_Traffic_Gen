`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
d/gChBcAYpAFcXOeHt91b46xtBsjSEfgRrubIpPCNWjZVn2QQYIoLoiBJ5lROjT2TFVr0mbEN0j/
51A105S+XuyGRj6zb+AsJQqRM36hYEoO/xyISbxHdrNAvS9FQVIt9F9yaT9vEIoHGfyqjDH0oavM
ssiKZOtSsSe4BbpLYz6nTeiweOmwwWhIGIV0oQ8zruJrtY4LbQY7owD9+R0Oo5tDy9R7RhgZUVA5
p8SF9ilJaAcHw5isJfCAmgP+kBCPqVG5jA+7IycfBmZWaSFgoQb3hhzb6b7/OasljP+ecggZvdGz
psSd/a3NxGdr5I9pAIh9yoKRgX+cUH9Z1lf+Eg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
laQzh/yt8VpjCEctZY2uX4lKhLuGxORtyEo0FnQPq7Qv6VFjzvo/kECz/qMLEqmYaEBHBJSVyIO4
/zzQPJF0jFpMyR8X4kCJFSDLPaB/rmazOoI6hTVpL8jpggVpNcQVfG0l9Earu1PJROITVIjRAM/q
YRUhvdBPg9OnFUL8hqTuKEqZn5quoWVCjuTKWW3EE9u1fJ4MSi5/yIktoSHpA7DktH5+78sNVQ5B
a9khdbIfAFcXvnGD6qnoP2Yit5s3KQxxZScbV/CNwuOYbiGtfjfuPYjE/Oiq9WWYAQ+TKqu6B+iD
DfqIfvR32JaUaSMd06HynoelRDFs6OOf9RY7vAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OEp/kY3McZSX6BQYBtRutZC60FL/ELNGF0zix/X/X9o4wKsrMosZC2d1mnRCl5KytKCMt2BPhYBV
c1P+BluvQA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CkNxNzbn03OcPbpELMYKhm/GyVj1oiKih6gVVaLaFRmvtexhDkHetzA/lxIYRwltT3yw3GJ5wy2O
Kl/O0ZbftxftLpS+zq2q2wDvGgoPo9NL34WE7LaCg/N6Il2WNCXe7weBKVfKG5K1S5rHWHn75Uq8
SJbH/z1MctDhr61oYlVLibn8DVMghc2DYiRfG7DS9N+NfmiJe0D4ya7AZz/7Pq40RYgNfEXSW6bz
XZUZw2vMv87xEPSbv5cyKXHfGo5jaPwSYlg+DevW97mJW7swrJzkGuId3PaT0iEQuHTLNO0K2MB2
s8nWzaX4l4+8fwYM08KshxHnemyheQlgpOxUNA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QjOidCUeKNwhQu2P1M/nalOnt91/DilHY3c9ALPdjL1tCCXX+XsGxiZUfQOaWTbGdmlnB26IUE1+
td+gHhjIiYAWigeoArqi4U/A3ltGlp6ecn6OLmakL4rvHmz3A6cXm8t2Mhlxq0aO5J0mbacB5wSe
2R/+iTHexeIaIqBnyJvyIr463If51nknVnd/J9o4PfkERDnMwIc7C52NysGuySRlA0dPoNX6PMa+
7K1By/gOY8He+Koz5HM+k0mijhOQO2P6gvd1KJrU/9KJjF5SkyDOh9I+TWwC78RwQWQdfBYL2J18
bcfUAFkh3XoGikaPtvJODU2z+KHaXHZXbiGwzg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
N9enhrcefX1tLMY0/2usctLLqr22Cwus4ZVzcQpZquo4yPohygb6MC2c/FM/HTONlKikW54/h5Um
/L8F0cFMSTtFAcKqvHHPZXxIloI+DFSVftfCiNSmqNOXVUXvM4dassRQo9kfNx8+a2Dv/dVATLqy
CTdINCYFGjp+ZlwtiIk=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kbaEymhSQtJbyCOLvrBVi9rdkt2DAELOFrQFtsslJ5az+lHBQL50p7GirzM3TBIX9rVjvEF9efW5
63kelPwdR0NLd9G2it/eaoog+bTByNZ8gnLy2uTr3MInvOTKN0a9VcFuCeRZ6wbnz283v7g0POWp
IgrsFEg41FL/46qnUn/cuZ77Ji9oEPcdH0abA1JG+9r0/1xuufET/SVlAXed+qTJyZjOVMUfFfUg
VXP6beh0mdLFJG90WXjwglp/dNhPvGRuLTfcfo7NTuovpKItqECJ1zxq9YPqcKQzVvSrrxYauVue
WyuhhuyjSyvUq3EiIO9Lg+X2MbQwGEcqPYnDCA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ycP/YbVd85MuHkzqUOhKjvDJsi0au8iD3+eblMS+aDM3nLS4yiWrvTB3na7hqM0purZGvgFQ+5Bi
xZqCj/smOFEjN0Zuvb7d+YlxZ0dCuDFipH2y1hxKv/YShodYIVy+4DTM3G8WQfNCuGsF7BxcL42L
qj5YhiWqBiwG6PhWKjMcLVlA1sLVHvra1fcH1xpKNFP2WFpe788qiOzIArhTd+9dTjVchpeHssCX
YwuDWXnrSYXlbXxUUf4vzzZr6D8uilDgWp6y9mEhTTpKAsi/PCTpOGVdOuSgUIsrLauemrauiwdv
fxy6Ift15ODo104vRcMaktyUWXBUKz0Zkkfg2w==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DlGk3sfE6Lm7cB0PQu78ecHVt/cR02FE/iGRUi4nX2ZraiVEI0WGbFLbypHwNkiO450wQy9eFpQ8
4/VVLYA7ZbviQHJsGEK01vRGYjTXEqZv4QdAWwsdGeeHEdm5vJbnbIkrccDCgHrYGg4ERoj+kS7P
l98HS3oIQSIuXywkVUg=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hn7XaJ++f0p87SdXn6hgLBjcZ+26Sm+Tw3tjInDu2fHj45yJfqEemHPEzXfZwCsQ4T3I4nfKkWAs
kpxKJnkivHSWh14IryoCx0df79XDQZ7GUm8685nQwbEY08ebCkB5Nqaq/gJKYZ0BfBaGiYhIzbN3
N3wRTXipDYFuw1KYrfrUBSWN1owhJKWj8NIye0WY0/jXbXK1/E7clmKuDEkSAl27R/4QHGzyLq0+
lPDbB6r5xdR5E8ij1s4XNdLYfnT/nyY3miOfruL9qw14DaHa2D7ZSyvg7FpCDA4A3GMuvFIaYghB
nf+lOdWWgMZfZg4gdjgh1FSGUg1dFROHnc5i/Q==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
wgTVdnaT/SBdcybR/I0ZSD05Z2ez8ncTnLgPIVgbYhNedBd9YfCTz9lrWUFTt9nNBi1Q2ow7LwPH
4ReGh4kZ5ydVVH63BgFfYQB4KN5Wyo2C2NDT1nAsy9qZKT+Vpi771/wuM/4lewTEBhKdOjMzHhzk
Cq/VLeuINatQ2oGwhA6rtbYymVN1ELPZtpOpNRxW/ktwyD4OBfb6oz7Kqfy1C9o7xk242tKw4yQ2
P8jCnZiNgYjHqi7rGOzvt4WhLNMl8IW/wMjLMCJMqso3tFY3jfL0T8H7Bs0+PnoJnjJd757fiNft
oUXLJbSGFm4JR6OjowBqykn0ElQQW+IZxkVXDrARZxvK9oCiIVzkHM7XepGIwnFZwQNvJMC85tGw
ba7UzLhB64dPHLhSQZmSh06unSSAQe11iHYu75jUMgZdLChnhBV+D9qESScUrGXkQelhK7H0e2w4
DZ75DOCiK0jPtW2vJDU3pwTl+ojjJ5bjbUnlRwYGKLNEIxOIsuhWSAaDdVj6CnqhTrKA1E6NPqwl
EELe3zq+eVFqsehKlbK8qr8NUPuGlKDj20Ib+rSD3a/gpTHFBwGCzSOH3qQhQnjUEUv9WHzf4scX
/m8xKSBl9hfzt7BwFgO2Ozsj5Lx/QzajmxhYPuH+jie6fRdo1Kii0ALr1HRiP2h+s6iIPvHrAzsk
dxbjEqUKzedFVd2PDxUG4Fy4g8A0FG+tTnXfSaWVlhktD/ALSiMMIoOJokcJSO4i0oPqAsjdpzGh
NOkyf3/9eTfnLyh+AetgvVRc1vFb5uErlFYIyzqRvp4QcsTHop+/0k65oq+mySIifz2wpeS74Flo
EBOhUTvd8y50VXROxhp/wOtGLCyt7D93gJIuoRlLvs9iBpm5N0GQUtaBR9h99t9qoNC8yaq09Esr
2n2ByYH7fGNKBjkvy2shmwo5dH9yxYrV5CxKqzkrIcokj6cwoDY9ByjO+3FIiPaFWNDhh6MM0Z/F
tfKuNJh1E6veNy4iwbQc75Q4UGzIwEuT9RxMZasemDVcnwkLHR/EfCIQ6L5tTSpuS4eEg41zJMBl
5d+4MY/gU3dGF3pwICySgW2ru1BYTIDeTEzm9JDBQHS1WnjFBwgdXrNbwtA99d9eCzfcQDXM1axh
nXNPi2AsXui6T2rv3DIN1xfed28GKLF6yUTiFQiOTblx9k2dR2A8f6dTfpdnfWiCNbgIDlRzxkQ0
tndqQSyWSd39P8+V14L3OKXVVsWBO9TUiTLPhha29aVm95zRrdLlUBvvTrdh5JwWzw7eR3GsEaiV
YHeh29qlzyiCs49ZtdkWzKJADXdO8tnkhja7o8ZeU7lLZxGBuD2ZTcwOHmNTLzAWbfeleSL33ALi
bclFWw+m3RJ0MoX5f3CT+J4zfUIRs+tfe9hmcHm6OwM+vttGNQXuNGMv2bU395O6pf3BT+AfiRFA
pKLhExIegacyOSZkpHtVi72AMlD0ynGX2Fwm8Kt0nGoQqFrxjxNu+ldspIQoxdw/8agFgzmCzlsG
eKZ9oXCxvGjbXwh2Xgwm7YfCssuhYXHDa/6/gueNkYoIwf+ELufBoG84nn5aX/49sJnGU1eJQWKL
XhnVAIZlTS5f/BJ+RzFQC9JGq4zfsiXCLzNkCDakNsaRfWUWO2ansbZGv+ey1N3GORqW9pHAUbPf
CRTZ4fJ1j0VCgFs9DIgIGQIMVGnb9C+ixnU8RryEQyeEW3CVDMOImJDiAwIoPIvE7oy2HMrwu8mP
dNSsFlWkKNfX9ufQsFCNdrToOECqmAbjHkwYSL+Lhb7+yLu4jzvVwmfb45KbNFRTrXxDhJFJLeCV
ZApt+ATQzC3u4CZXg9mqneyaiCE+6LcCM6nliRTSJmeabEXQMMtInrtMWvDs270PiA3tC3nERdi4
Y2kn1ViyeOgbth5FLPAAA/qlDEeXVxYzkuMCG3jtU1vOnTFZJJYIcJ7OjF0sSuv9DWwm/xGj4xhG
JiGeMLZDhkiK3Gn9bgNtKlXi9HmySKAn3xoF5MSwgaoX5/ZZNJJjAFTaAccVceg3mpsLK0VPU76v
6h7KAlqRORp1dUP/eRDrGCpUenKXXjW09g3Z1MPxXJ7Yji+TvSZZ3PlYBGY1EadMnM328dt8zlDC
KMvQtpUVcH60uxnPjCAeoGyA5NUvAR7UqWtmRURfKT4pl1q0rAnNnZhQ43aeyhZq2D+RTFTzTH7i
uQGi4Oc3Jg7eTJQQoKd6UFz4UXPAQS0YlTC35U5kwmo2x0XQRbtBW+etz6h+l3mp90M827xm0Snm
WDVbkaustCwbE/nWfWFMC5HnRargwnfTjI83VGFZniHdOJLViFrh0fdHS/s4THRUGkjAi4IzFkUo
HqHNLgHgqpF34V5CeT7zzQV3dNIhodIm/72wA7r/0ROmhElu3KvPir92NS5F5fx7qZgI0EWuyDCd
DU+gnUQdOlgyiODTZe//pZ2jsp2X43VOe24bNAFPEG2SxsebIUpVrUkLsytWmX0Zu1XnNlMP6nsX
VmRXskNydf1uEAS+42yQn1cYstGecmVctpCn6j2fufLtAo6qgGDdJbx4z1Sw9yKylsh5EUhz7XLO
Sxl+s5YkqVqHfeFibmQQ76WqywXLmvCKVq9QgTf4SfcB+qltsnG3nM5Q8ignNiBKG/2jKqVcpOrH
r1JBsj0gtXDhuZU6l5zK405UjiegX6aezUL2a1CIU1EqYaIAmAleAzrXbVCMJ5Gu4SlrRsxxA/0B
OHJeH7AePl6OH43OfPXV9yIVSXJldYDW+1gM+7HlEmSLYcPetpKrItEri9sVL1WEF7a/pXZfWeYQ
+Q7xc6tgSWGlrxQPZYd6Mjv68kYMW7bjM2jhWdF95rzjfFZbj+A2DyLnAVZMPng8Y2jVPvKd1M1s
4xs/M8qvdAA9eBUL2Ns+4o9SGxWvHzaN+Vw/Mrctnm9UPnTVBcmIP/lN1kk9XwXW9tEoJFOzt7MT
UkfXcSEmW7edRr9Hwb1RhkTiOp8Aocx8vm1sKVmv5fOZZVPgb94BrZpXk4MOQ7/T6QL7uMLSvh5A
aNcQ70SvOvV2rn7L7i28U+gkruajIQ5+gtkicAfwliYtSKeS8C7g60fSxZdThuHzb1LpBFWr+OF5
EmFsPGvC85bYirKib59N4IG3d8kpIPoXss7aseRoYiLXqkkGiOqogpkpltYuMxayngWbwzwySbnU
3TJ03IRjjDevm6NBH8bGLYmz/f+tOxTBfWssX9Gqf7elDZZOstBLOwuYOkQVGahOmF/Gq0Bt7Xnp
Nr4XBcWaCzD1fLfpO1sdow5vyEWv0ql2KCECR/fTI6eEgjSvdbasVvujZ/3rFQuIH1a3sAfLcIt5
tbtP3hv5uKQ0/eShk4NxELz3/o/y6LCdqLcRDVK0B1S+h69VdRpe5Z/JH1XD1xFq9omxQ4jzcaBv
ZZKaqosMeh5UeG6GDvwZN7n6l2N/Ee7MNKfkPDulLsyEE9IbKkuynAMlD/8paE3HLNVioUqt3I73
x3wgq9yxtCAqFKiMt9qJ3A5yfHtKRkeXMxsD/OPAoUJpoxSLaatUIJs3m4LqtdAL+RV4m7qQBnaE
rLYKj2kmDvxQpj+MX4E/PqQtZ7JM25JzE240dQWK7sGVIaa3kPq3EWPuNQo30lhNDdQPNNigvjSS
ZEP1ircqKdA+QyTH0cYKLuK9oEPy3Ck1xA6J/plsd1lIU02xfGEjJa/f3DlZWtnv2skXubDL4Obo
+zMbd6sxML3BBT77ao6yswZJbXt+JJ38mIRRrRTrmdrpJsp7CnU2L9oZU/doUarRWqF1ZaSFT3YS
5+rQkXOA1BxsLtjv0q6QSC2iMsu1eJvVY7Wp/8EAItNsZ0XupG14skcFwfZLjtRpsPwDxf+w85cf
CejQUqf4S4v+t+W98+MAnl1Wkj18YMaBCJb/D4UHWGhImcYnQpUYb2FmkPRTcN3+Vhi9UGeds4xq
/+y9r9kWSIUCZw5DUXe5kRUAA6E6KZP+ZACQB3w8Cy7nM6wts+j+CuAgMq4c3eDv9pOcF9bL/oW7
Xq/q9MnhJDpaiR3UYuOa7sd3lqBUw5RqrCH9OLpn8lGpnkJeC9wqMZd5Z6OLM+l/zv8VfXLa6inS
LVjivPNoD71p/z6qbU4QRvBR8xPx74PAtOUwPqNXsb0Gl8p88JNs8HWRo2iv+W8RJogInvmHF6c7
w8BYFOryEJLZ9npGAwRGrVza5ruzTRaxQ5LZkkDLeW0mRktq2u3HZsLLgZZ0C2duajs2fkhhZg3m
538UYqQD97KHPAnCT7f4q6I0z0VhFJjOd3sYOgQglJLgRkrfgn3Xn0/guMMqYKu+2jwe82cMAV7f
wyTBd09MOyEI037Pblx/nbkECjzEER3Wr+vsSEXGTBUII2QMRxLVDrjgn2a/ZVaf8J/lvXY7LW0T
qq1QOHnK7dcSqMstqboLKgGn5XLpwSiT2oQqiTf0JQpPj4b80qp3CkGLy894v4r8hgm9wbKdg/bH
/4L16r1I2FdgpL7yeU8f1uZs/+MjVaTEXh1aY0tkegzX7mXstdDKtLF6dV/8CSwO+M/e7YXqdfd9
EZ5wqnT0piuIkiEloq2ou2u2TZRXiQyOk5F3GtPaINvwBH8Uc3zFgyvpO9syxVu9wo15vceoxX10
RjnfpWSXfRb9CsiF0VS3YuudqAyfDgDfZi4yrwY35O+0b8EpfiqdQ//zk2zyPb/qz/eH4/iWvEtR
Rd49d7rXW6s0q+8OMahbQnDupw66myYOez8HTBQ7Hix9FOV9HAfpYXhxKtqROWlemF9pa59GsXGG
yc7O6ZUYCalut3hch82Ch+Oqg/tCH2/f1W8f3GfhQ7jX5s6N+6H1MjcTVVKCEEoaAi4dR0YjZ/sZ
LchPPJcBLGGIjB1aP9/vL4B5HazAJpaUDECPr8e0SZDJv+Ty+zWeK/eFEfjF/y3JiMch4lVkgeMt
fG/Wfx2idZyonTBSLZtEzvNTwDrIIy8yTNEuFjE6cpDsprwe/iL956+pV6x5J3lg5FTS3SnEaZKI
5TtCdYIAnDs0BJG61c4bzSCLYxRzx8K5DbttTZNBZfne1PLIBKIVU4GLjXfO4M/lo0LJwd/Ylxpa
a9jGQQHip2fZH1CfGFqTtUATdgTOWr2P4qDTzl3GEEPyFlDTKYRC25Y9jpiDKqar89epyyzjXGFl
ftL7rL2XVUCko2Oclo9l7hIPVJrr2jm+OApSPWhh5BvjGgzseidZjuNsmZyTeEsmkWYaBF+QktjB
D7eVoZIygIxSdaMXVxS63aVT/Vc569kr+cKAUxlFfbnN8aO1RLEMbzZMFUhMkxM/8lPLe6LyqVik
3GZGXIsJ+nETSR+sJBHLi4h043+nO31T6SdjVGxXOnZT32soNytEuefBA+ckFc6nKPgC2mW9KRG1
Uy7ZR3FPm1005OPJviEMjCtc0BUEZe9Us5d04OWd/jWms0EfaxDYJZFW+72pI+1DqWFK53fLJUAS
vHABoA0J4DshYem2U4LkOUSB3vlENi8VBb4mh6YXLex8P+Eqs0U17lEeukUEZunTWH+NHLYDKOIz
09rRmkFd0lnc8K5sWx8bf5d65+syyzwESlYeOM5T1lFuLYXWzv59zyqiAN3DkWI/Nr3dZFKFxCgw
KK2BkYfZHPB2UmVIhPE90UCsw1vXgALv7So2lK7Ddhy4uhBeIeaEADVXFCr1RVj+hTopjvCCNXiy
YWWUrM6ySJ46hotxBiOI7EWFSWMG7ldQ9R/Ie5IJkadsbxDZppgbg1n2OrR2WcM4DdI8qt8iQX/U
PFPAr42B7MpP5oWWy9Gd20zoiWyAmGjQR4yyOotTep47x1Juu9uvNu6IYFvSJ9IUmnxVj269920O
Vs+eu0HIuHFiu/3MvowifhYuLDauL3iWCZ+fyV1lws54prgSPPE1pJUmYQMy4NEvAfYwe3Dl/j1X
aE9jtuIutcHUsVFTG3aJKlbnYOqY2FKAwda5SB0eyOB43j/9sYk2sqBsOy0ya3SuEMTEO6+vNCIg
RrQGCqOr3Q8yjtT0GM9XEIWPgXv8RuDzZG8Hrn1TQl4EDsJg+0XRHnrob2BraIHCbrUv5OWqqr1e
LcWJ4dGZv+zJvn4nnHbEbOVt22+khg8TJx75Hctj/gdkQ/rGy9x0KJi0FD8/jG69K08kmXnpyBxf
POPKVCTx8ut5ZMEgcmNqxjzExb6vsuokMQBYF01AzKkIm5NsXkBmdxGl3QWoIRHx8qL6Kz/Lfl4B
KyPOkFlUw0nlJ/Vr4wloTMJJSiFYFSX3gH3NBcLfkb/jGXBRUywp4091uIw+lAAA1rx3ZemHJbb2
RtOxIZ7dDfCMsUX2l9fTZhJUT1wFKLNNGlTSXwP9JpjtW4O4cxpCBXQK+QXe9sq01KCVv9t9seHz
KAsstyIcO2PKA7++A0FQAwg2IBWcGlz9zSV4b792OxcQxXp0KexwOHsd/0lEqfi6bNw3ihGGSCVB
nv9qUnP/l9HqoT8qfzq9TapRHWQAps//SJlm7e5EQwEjeTfJv5ZeHfz5hH+8uhrAzJ4HgW50ko5B
wtxYRBDrW50MjB8M+3TJ2RQY/A20hi4NYZObesVz8WpSuvmq/6LLAJ3Fo6/bW1Jy3MLeDitzgIiS
KclOGGRwANbqTDOwVtymQYxl93/rpqhRUXg9tZI8wlGvCn+FAfBP9AGOO/I9PiWq2qA8xp0tlMrQ
cwMvmnam0XTmDGdhLp2QKdle1TwliEU33HjrW9T07mnaojynxJ2x3Uhc5+w+W8iE+nzZMmvyuZLW
l57+/xQDvHIzxL5BcfQ8Kw9ktvHD4+HpprgRjopTIyeEAPibzkxiDtQvf96KPhBfg0gfsppOH7MQ
nGmrhSUEgCQEVKT4LK6O/3X6FPkPWGHBFdLTti6FIw7onnjdVFsi9CwiNo8NwxhpJovMEhH0Cm78
XT7xvUYSAPW2ilLqqByYNqlDbwBt9OXSmOkzkARivId9bOI/1olQYc26TmSMXlgnYuamoe8kWUza
Eoeg/8J2yGOBtRMPp5PWc6p7O9KqY6NCmimfqxXz+xmnj0o7bgnh9AkTPhNZxe4drsliFowaot56
VqbT4NCnvOIyDQD9hdq4qHsnjQnJlWPbfe3nGRsDh+hQo2cQwkYT8Hm0b2kLjgGgliHrZUpTk0gU
O18UUKaQGIbJ8F6kVH+C3JxjjRWjToneIHasfWWMdR8yJ2Nzk49pqwW0HMTHKncRKn+8JVPZZBTZ
YFWl5ciqISWe6sF0OAQR7xP/Et1Gmjmt91QZ/U9idxi+eUFo+mhOlH24dZRji6ZIXoSP6thx1aSs
4MPOfMvl0uJGvGE0M5QyOBW2eD8vLmQOG6u7y+3ctP2vd5Xa8bvu8zOYSJgeKHCSr19x2H7e1gbn
5HD0VZx4t/QuFdI6893SLWw0cWSgccwvCc39oqzvP620HryZqbC31ZHU541mUzg5XJo3qce5BRju
RZcoDB2ka33uCofMWGRXN9YU0WTqhHNCEw3FMiOR1O9JQvtbsZbUkMaN2VHsIETS/9OTfhhy378d
nfDgOLNdxUJnylNnyj2FOgN8x8DLA7v8TnqnG7OH0Y4vJ2ufOgJjXlC69sGNOPnn0zUpxVs1zVXy
5BoWCsXREhGvf3Ky+aJZ9GPyQIpwQ5/cH+D7d5353JGXoYCfRXRPlJK8pkbtvsH74Dh5Z3+oge9Q
TRzJMDuAZaa3a4DnXh6FDDna6NEdfm+GUOvN35Qbz2v7iG8lIZzA4k4djAmR566cAhqM1XyzNL9G
EvkYGBt8plXqD3cEtx/CDCfnJUcv7CR+Fog1F1WlbNH6Deqjtyo8k5eOySqJKICzO1x9lbQZjfwj
bIBfEGolniEgk28NrjlfwR62uDcTRjYZbmKa8r9a1ftDsw8cOWDfilHH9cvueFp/mMFfFI2zVnRK
W40LuiV/OXdP+fAoMvo0TmSmG0GiYYt4xa6n9r5EjgXlJpWsD9rIyAzAHW//powI/lYBP2ayUwyF
1O0HIPzaclNZ3/3/18L652k3ZuUlMlNWUAl7IdnF9IPcImWy40v6ZPzyzID7hdO1Dalhb/hN1IJA
cITf+1WWdcfiAvBbhR5epKuHeCjUVaJ70uhdDZheXfRTKKe3eqK7KS3pK7COIFrTawQw9I4GBI1w
UDADNPquo0XTb4dklBkPmiDFsB+6Fp+XdF/zNz0nB/qnGE+rtRMV0ocqtjfNhfa2Me/0B370KL9J
Qbw7wpiEU+HA7v0WxdeZWtChPhyAJXwjMalGk9gSIZwvR17SU7gDPN4H57xfClN5l0gkkvoOs6Qw
DF7BZ0nrJe4I/E8zJoZgGQGEK2eeiOwBFPuTxrZt20OS0L5f0BcNey5LKuYqsCpo4gOG/YACEAA/
QoW4EP7aKYgN5uB8RLdBSWczxiExcQyt10VjKQJkYh1f/ZvgnpzJ7VYIapBDblSgZLEEefP3SW9Z
VizX3q6tjbMTCudEbmbOu9Nw29a4jr5LWB3+6y4SaGICqupgm5OigLQmhSX+44ZE1nrjTWMWPz+Q
N2+fuHX39htSxFBN5OqRrMTyBK4/oAU3LS1mmVHq99XU3jOUINFxL7YQ/av+8wJo6/ms1zB4z4zh
XtYvnzg/vWeulfzbLcOjxUceQjD7XQ0OfpQV8xoWeMUZTIYArT5Z0d1UGmyrpjQOm8Vcnm9dj6yv
ZxgJ2D9eqBFE+bGRfIjXyJ7NxT1IQHZhUzcX8YsaT9xS+vV1ElHHsiTWHcZ5F3jC4TsiDIhBvnZi
QJ+LrGfmBt37pgN2NUt/VC+OAPDDZgqIflG+KtKkf95Cvbhs+GpMsI4jOghX/sp3faMSWMKgs0hI
M/dMrtec1/96km0Trh/Cv5aholFJ8nL1Vdn1dftqsjsFUcEHbTjYfbixKFRHIwDu0tWiNf40+PNo
ZUeJgxP8llH5YQ1dra/Kv9bvzUd0zVaN+lBEvA+vBM/txc2jYUfEapXdbGLYh+7lRY++PWfyFWrg
y2W0YJW26vnb2dBBDU3HRbE5cCT/wnmDmaMBAMW7CHOxLGxPjCY0QkjDW0jBvzpgtp6pw+tGkAOC
A/s5balyp3XP5wXmJymPlRkyXJuOuq5UyI/c47Ej6/wEHvk04LPU91JIwmX92nCLddt7iHR8vGjP
LYPkv547XMBFSxQiw2l/UjeA1DTEUgorE89oJYr8wXwjkvLOI+p9g5L2aiglDdTZj3ouqyYqV2r6
iMDR9ofyk6JXnuNwEvHz5fqLN4za1FJipN1C/eOzh8GgmCMXYxKf4QTfE2qT3dVohanNbunrS+Bi
jWmY+UKVfqiPEZFCxdsSeYVNncKif0cyvDVgEkyPiCGjCXv33vz55aORrhLbxXhrOVxGESpk3Rg+
b1z6doWux55VSZDR6YTOC3X1KinaMo3hmGFsWtj6AOx5pf+U/xvAQcVUKTKWN1MPAC2L5ICFK7HB
mDdxAys0ClvKikKDb2CaRfTWmslHXcz6NdQdWKU0ZMMwhcmRgX3MshOex1Tnxu7XhVWR23NwClhm
eAJT5dv0/h/QK9ih49KphDWzL2YwfUZhym64plD9eibhDK8zemcxBjfsGQpuVHxlKJ5B9p3hhEFT
BKpeVd1LSg4/QTp9ktlHsa9TR1guiVAwcV1mUB5k8jkRPELIjk7Qve9Inj1iJDHxKiDVfAtjXEGn
SbUgpyFVuNq+Dxby9lYOAsUpBAzk8q+qffp7jQ/JYkUXOrjkME7FuARa0W2YIoOwo3o019sBocdj
F7PRhIMmpSrNdCrqAKKRjsEvt6N3bMOrPnFvxOtmtZny1yCNzEPOvtKaKtHDB0CcAWhmnVK1Jw9Z
DJWk3WBjwKh2YEWrZzWnohHyS7wuezMF65DGSyGInErfLLvKWDqj+ebIFjfacQUS4Lkiqy3BnwbN
CELJ7GTQTrsiF9H1FycKz+rAbfIW4D88qG35aMfgafMvwNGRAddvspvXWahn0DkQch1UjYK3MKk+
FJUurGo4WwFm7hOwW/+Mb5Hk0+YCOxKnWDt+dq4DeRKbfh8jIkFcyOlg0dafeS3fSVSxomWEwUFM
72Bh4GyFjTk4boeiUPG2XwVE/AKUZJ5SXpls5DRu+8V53s79EM07oKbN1iX4+1wLk95nsqs0Llgf
tOF4DeKiectncHzj5v928rYxqBvdBRYsh3xeEtQQ1q9vQ3hbWv+Vf5+NT6XVginh3CWos9kKmmMq
wt2X20ieHJxC6RpnkcqfuhLgtbp0GdAfxwXSCGJN77nNWX0U3FobpPrAa5WCHD/FVPxhgIGYAe4j
xsX7nSw6+yBXA+YT1G1qZAEFtA2lr+FpdL1lf8Ec7quJAFdrJ35yZJC732LJEJQkw1+jI6MNR8en
q6ivj1eGLrTJYe3wYG6pAnhJScbKdMEKOaCWmfpe2lyoIfhQuqRi7Cw0NdQ5WLED648PL3cpsNjX
Udyb2hFQesV4tKZLA77h4xZkC4bxf7CZ6GTqVBaIX3eSxkeR66cMMGsN7iz2mlcGLtE/Axm+uFk3
5sWeK2GT/lXweti1+/HD7Se2i+3LMcgyhr4tr690Q3SWIlAn91Pjj/PeIXwC5Nz8hFrNRzs0GvJb
RqwDSPn/nnoY8LSEo508PXQtyHewZ1isjgyEfZgSyL30P5OkBAEzBcfCzqmA08gdCxYA21t0Hrgl
sFB0DdcvkempxMv9UlEeYKPspbtx5RHb3IAdk+vF+SXkdvRGWrSyjMxHfBKHGB5UrYbefhcHzXmz
sjiXC2q/DIg6CClKcY1PqyiLWeGxhRC3bNPRNKM465fdqGgpDYFGbIEjWc/Bf6Dz4YxT2q18VnOR
QryaeISRhe0rLGPmuW/1IzuYgeWo1Ibb9pdHBhERoO66XokWi3dyOjghmC1c/ZAe84PBtX5ER5h1
xbShRu/KpEsK4lbscRu83gtRb4MBDaZBUFJkfe/hC/5m2/k3qL2GL2MN9S231chnmJWtwC94+09G
OxisCf0KSnU63//+Z/seJ0BzAfEnxKQM9Q06Zx6e2H8f7D6mPo9Rx8/rpi8k7Ou3leL4/QxHbXHQ
eXNbDSJ8ntqSMToatbEPzEUay6bgO8SqZoiNS/oB1ho/OIJwxdxgrr7T7YPvVJIm2ALuT9AD5iLq
OOOeR1aEwLyh5nbUnGVbZXrk7AS3T4vkVHDm6oLXvfYDu+QBAuLIXepd7ea9lWTaBA8QrdPnJWnD
mhPkxsub4Cop/ajt65V85J7nvZPCpJzgXFshrFzd44zAtbaCfA+Pwx2P49ZprOhACUJaErAJhoGk
HwaQ6CbepTDJmOa1K4Gc9yfcBwna51hnApVvGK+qg0cy3hgaJ4wFrEJvgLsou8bXolPQHyzVqBU/
xnXM/acedn3Zf4zULKviXt0CTf0penB4jjDbNwBgLXRtekxJoDt1LLbN1/uQB9RRSPyTV/3CZhPn
c2ULRk4gtBS6u0fPxyIIryuCdtq61BXOESEX7pWvhzu7LQWaQoZnAwzt9zBHnHHHj5O4D7MiimKq
CwggNv5RkTcrVGkZdzcVOVCrRDizLt6lJBmgxWbe0liutx08SZs0VcQQyviapSqDELjuJlLWtUap
Lzvrk2zKWe7BEOFd1N9g5mww+MF3Hq1bveuG2+w5XRYjx/Oa2Y7oK+cn+fJ85hD8U1mZa5aspta7
hSpb+39oZIAqVfrcDJ92lHoK15RFwuA0a8xfHW+7VwnGi9cXMbV1UBAuzxeuu+KCwSR3K1Psl7ve
Oo+KR/eCVWdmL9DdVRpwBzplSSXdeI2daukiwBEcz+ZaW8ZAXh2Ov258uNy1b9GBc/VzfRcx84am
OEbj8sbHvcUtUYNmt8J6/M++dow4+ZIOXojr+2APnPjyHi177c0xRnMqTGvVlpYOBdsm7nWWUvnz
eTGlnEoNmL7F5vRD1G+gur4K8AMMVte4gF7d+1TMOJm0jArNGD4XM6OZdBtaHDfON5jk3vlYod51
JeTfSk81hzClDEYBtTTOpJoORS8AoCf/hRunzuwx9y3y054e369cxMKrXWDK/sFJuCZ4U5+2Rh8Q
6w301fUN9APqdFJuAEenDtPGfqybtNuk3LHZ7z4PReMO8H8KKD4p+sMyLrKOJNQrogQ06D3CP+xX
M1CbsubBSaGmSJyKvo+SUfwleMSsPX2hhx97Mxr3VcMP6BJMQ0oJFfXPCu3MyqDMzACGl7Mq5ojP
vRvDV2vsSDBKejfPQISEN17Dc6ro2mpgWR0yjGV9UYNic/5RZsK68iNF+E7IHNly00gD1+Le0miN
YiXh7xCb2Bw2wsUupbvmhf7ejTtApEDxGdFeUQX8bsP/EcxwABdxw4sCl0Nf6OsWTRe2SIKRPiPX
G8HptDbmfwtzSovfLdElRdhetSFQ4T9bYaGt4ocYO9o2da3csIl1fROeNSRnBRhTU/jxvYq1KTCX
L1zBC4WDUkorPjtcMfxnkQn5MofBJL8HFn4gexsQDnS2qRL1U7g2B8Ehc12uusLEHraD2+MaCVPr
frPNKL6L3GbeQb/5C8uyCYXMtFvxvXZV+khyqYKprOPUEj8Dhxt+5PGeyGrH1g/A/EiDAXeEj30i
PKwu4x4Rk6/S4ThfyivpjORTDU44zQTdtQEwCwExu0L7iddvYRAtVidJ85rUKw4X56Qjc5IbU8wS
QeOP3SmFk8CTN8vtbvxGRQdaE9mVCG1WZqgomojBU8cEMLEe0dIW89T58Kw555oyYh5lzwjOJols
Qdm+YHJ7I8Zk1SbLkUZjEPka9XlXYI9rYpTuJPMh3izn0ow77QO5FvGQ8gD/mbiuc7+8GMDVvY3v
NzjkMDNrQ5t2tJcB251ZK8Kic/bLADV7C0CAN31AGqRAVsxPEsXaFtZzyWTc9a2Kv/6dOLDlNBCv
LUcoOLqNKZ8mDGHPFUTK335pApqWCKRgT4wW31SvjN1IWCGVax2AZ0hspaEpVpiAtDufgbCcMSeD
wW5znzvYOEivS679siJaiBBYwu0caZwujE/n9ToWN0MzUSelybTld2Gl7qx2M+wDiFT3SGOL6Qvk
G/wTpOApWYkrU5ypXgow80L6VzE2Bec+moNlmhuNB3SbE+CK//YtwdjWD4RvwI1dTwuaswNPuCDV
MpQyBmd0xxH8BKtmdxFSYj4okLED9Okc/5iVLYMuvP7HuxXHQxBxAmTcyi3dEmf4AHWdbe0o1KgK
xqfZTjxehsnMDCT5xLBdk2tpIS2s+HLWTqu8/kifrst/DojzV8nzdeg1ZKv+yWKfgujiZv+RNzIH
HRrF3dJ6aZ2Xrm46eNfsS9jMf7QKHuG9Urk5o94XskVAmqXXBuAIHW1J8UtTK75dqUaQ3lrSCjy0
YLDFpuGRqPCq9n1SV5q0Rma6BsUTjgYwtFKeb3o+jRjwSaG02k0kxVj87OALE0oAa63MVN/Fv+p+
pMx3kZ3piHBDWMcAXFUQR4+UklpE51XVZF29WTn8plwdTgcfhjt9OJyt1QBTMJaOs8xA42b2bO1/
qATp0YdHcykj2wbi/a5EaEaPMygt73XngmCis3he3atK0FZsHSeZ6lkwQXHv+ULp+mzjYAG18Hqk
ovfd2FvSgwEI6Ldn+3FD6oSD9NMNNnIjJPL44aub6Ku4EPrfNLvLF0IhidBndcJZUxFAzvF4s6i9
Zr7tXVr2azZdKwB54Ov0px5u+lqn0MTp1Gz8k8xmH7fAsqloVq5OdZsinYRmoc4pcIGtKw3/i/gc
W/oVDoTS6mElFfgp3dknvxp4bHEPK05DO6wof1aOOLHZok8oarm83RWpL4thyD6byi8P1PorqZX4
SC4xxfN60j1ps4A9ruM9DZuPjujt2FRGulp6eBAcsLw6NN3bFaCQbJDtlw2EZCpBUi0kXi2nca94
Lx6cq8x/rwvm/dz/hYrT9vSYsOjWgBG6CV02oSjy0n5itKEUgtVOhC/KjzHVrfgZYvERzm4YOGEn
Sf7rJx3rcBgQOI6hufOP1AMC+7DRDQ1fQxa2z+NPtOJ7zD3KslXGmrsP/MdjGxQZQbzR4MtY319s
SaPd+/K+xZs15vjVhht0yU/zU8lVJbunDEwbRobrAg2cqdGbeGa1Vmhm+lC4kAUGvF3z0EGG8HtL
eD+g0S2lhdg5DECwKev9/Ca8LCR70oNJX21AnoXYrha7u2FZ0Z2NTHUv5qCyM0XfH5H0f1EU1v4A
yv6RyglKIUewPYHWSHbkeUODI/ZXqhK7fBZyKSBv13xJmkrKhTEACWIvl+QvCrA7IU4UGrrtTnjf
ibePdWHL0ybGNTWivs46Y4nDlhvWDEhqrUyS5lYRg2I8+N5Pzbxm6ULuJQZdElt9WRKrXsxJ7uil
xEJn3UNBWQNLTW8WNJ1hkYTeCw/CYQfAo5YAFoH7BOQYPpPKg1h+otoDMTpHWASwmGNgQYoe1Ga/
MWKOQaC29yNc5EyoZ3G622HC8bHBw1FtWtPaGDe5LYLK8MzAPwskq36rpYNW6iUb9j7iZNePuWpV
BlByK6ikKVOyylgI5VTZbrkwGZ/eK7VwzkTON8O6X3cTdLf5n74joKcCyeXSg3htY/aR1xcN6+0u
7e3wgce/tYadJpmtkgEtrOMZrW+Xp45YY2SoV0Bhp0R7U6JcnoZJkqWqCM10Ci9fOf7DkjOTrmPX
b/EsPCrqAiH5SOv9UmTZZFrGm6eTQ/PnGtNGGL18d3Pb84aRh9DJT3c0lPmkCYKix2/v2EscIdBe
6XvX8CX7rF0Plr9d848m/UYBmqJOQNPkKyLByz5itWGzdwsfHJXz9FOqveFRPqqDSNj6fybmzhRP
AK3QIW5Cec07MYwxyx3w0FmIcnPcpiDQWFqhYqgYiLKZQW78xKuideddAVtpUaeB5RiXUCHRcUlb
4+K6WHGpBscaTaaaBL9KCJ/ksrSvD3k7nFGcPW9FKoKLjGgtqeZDlVpqeyzdFewASp4Z4v2EVRAX
qF+Tm8ZWqTImhlF48jROhqJ8k5WcN6qXtUK4LA1tXEd5xITUsFjw4KhhHYc0IWMXFQSEglpL372A
huo7KZGeVUKAanWwvx8DDnb+XtUH9LM/IudE+RrHa1PatAjpruTJ+jwopTEFjPAYBJuJ8CUXz3uf
gYFTU0K2NQ7hTj/ksBPq9x35YHt1zXNOW4AC+CCG7whTOPaRcjMnU/ipPiWfZ88aUgV8GMydaFPo
05tolmydQ/85+iaZKg9H+xQB7nq5E5ZUEWc6LOhEs1d5Uu9svWTHZ8IfuPB/cZ5psEohS/rY3iYz
dCA5nL1monA9AyaNSiijKbHxiAbtXsfmdRTI8mXtIzU+ZfypNJiz1H3uvEzMtMKBSlU+/YFZIhui
A7bS1LBLS9rDRIa2zOPDzgMTygnf1SK/MsDw46Xd9luSu8ksnuuBTUxTq0bz9Fripte9sLJkQXcV
P9t73HwzjB9quSvsrGOhhKiMJWit0oTqmgDI/ZFJ+CZDSX824t+SkdIhzHrLtVelGtPXyrCBX356
Hqj2NFPLIJvAsXXpfUtQn3bAS5uh/7hIn/wrBOnJ08il/THpEAvg732ZOc+zU4xuVISVrhE3Ovg6
V18NCVlX9UKwMcEDFhQws9p7dcIYAB+2/cxKYxB2t5mFJTZYTi4njmDS76yBA2JlG+L4ZydJqj7O
lb5+/QJEXwF1p7jSaJ1DT30RA7IKmrYFt+E4JIUYYBZwZKe2m3Ouw1nr24j9f4eFzpS7hMV39FC1
ajfjr1SiPAl6UNM3rnuVW68pNFu5RP06XFGaA4TmVntpqEWlXly0B+uoo2urCGXPsK0Ia7jVYrF+
wiyEpEVH8juEbUXj3xHXzxzHX0zX1B0SKp5Ihe3DXEPX5P9PYskrBpHbMZHQklKNO/UAiifx/tQd
P90fgpvEgRX12l/3Bn8AYQKsXC/1qwuQmRUxyJ2uhrrb6l8a4EBOIQduVK+6Wf4I0uEWOQOzXMH5
YTMBsSqs4xGkE71LBm0gcqyUt6DvLzeJORFvsU/7F6qw/S4zojQ1QX1WBm+2Oykxz7+z3jp0Y7ls
9nNYYhtfkB6dfCSgRtRFlkUncm9pWt/glUQtieOLmNJhk+GggoU4haIfgIRQKl+2opgmJy7Pgcyo
WuR0R9uH80zbP0Y2b6LItFShUiNAmGX+HdoxY263Lve5FGvKpVd3jDCwUjLLTt99y1Qtgo8j2YFF
OBG5o9NxW/FUiq5zTmwLBx6S1b5Vfz8XjADrJks42CIKlvd4Hln0E0k8M/FyZjE3YX+ml9qUFi7X
PEv0v9u8Sgj2+g8r2CyW24wWX/GA9lvz5sPOljUPrLv7HukUE7zRtUiNoowouVGo167Npnh6RkSL
UJNa6vG3Z1AUKpXMvfSBHFAXJ0v5aUqQ1Ita3bEC+WE69wZMd4EML+o5j5Jahf168y3ws21Xi9sh
bARUn0gQdghvayINJ1LqFb/A+j4q6PDkkkR5JeRKsRkHo2gB4qoijSSlQOU76QVAeX64swnw98WA
HYPpwSIe/oTA2b2kMu0IL1SFiZg+gH3BLaiP3HwBfoFHYFinQx627FESE/BToMStRCtnTuV3dXok
lPKlJMO5AfI2D1OK32Ce57H3qn1qoSs4tU/DfQfK1aRVcbO91gDuvfoBjjsxySEkPmAyb6gfmH6l
i0hPf7QjZc3s/XgBuHm79ehnApkZV4EaPbAHzLeOYJn+8gSeusPdTuYphX/fTVRX1xbTsgmTgujo
YlClK6x2sRAwPYFF/xxYcJE8QawKMHT1K16AMg11AKgaBatKTWf+UdW6sstJ4/bUEFU7vCpj9bA2
pIpfs8fBuKQLVhG0IA4E1IjNaitkP+0XsU+caUfs29gShU4yCjYGgb0YnRxahEprV987GNaoWVF5
9doeXCJN70m/Ox9eVcbHUliJPDZEZ4mCJqlSd5MFFGPVo8z5jJso7ha1aSsqUC2LW9iznIqGMT80
WI8cZRdSq1V5tW3zrlR+bL2spQQ2qEYfB7eLafNtHudwqxxUpqn6yskiHPWuiCjmQG1UnQvpN39M
aKxaHC35FaYSTp5M+wPdFANobDLV1MHMtCkaO4yE426Bg07PKe/aceJJb3ciiASRPX5Jpet0dPn+
RrjBepzUq98owyVW9HZsdKgkq/ibC+Rw2lEt5qbTOa4pP6kobBcSFh+a6/ofm7AIwUSKhOuK6kp5
JSs6/oe/PjTxsJe0B8eHTJVLueOL4kz7/3rcca7YEqM63IS82HMmsJVI83CIw2onupd4u30p6mXo
uWT+WIjAZQugoT3LgGMsc2KX2kGlz4IXXc9z+kraNQUFPHFDvl4+9zH0hPm+LCP9E76kRpcxEFVz
lTBzL9Q1e7Vq02NH+WcEVp7PS4VdleCm3QutJJMFJ4QVAu6wzC8Cp1SWgrzIRwSwdKMxaVLecDSR
a5NXAQYUKqYGoDoU6OURJ2Q9MDMP9Wk2ccdr6vrQkBm4ZJBi9MI/LEUGYXh85QEW3E2hx5tsfug/
mxaDeBio4lc5jGEfvLCSPVrpwSUN3+kj+0+7i333rMQUT509NMpnfEQuCiuOvom6IkRek6hBHZHY
jtpScRrsejp3uU7e0yNr+SYBBBct8L85NydPSC5QNqvst8Z5/KG/lq8OvMrY/2V5Wsx3htQ6yO1G
xMeY1Sh9i9cgvxd/BAvR5iLWMhsovKnCcFS/gbmtLtATXcJi7G1mGXUO8+Noz0gsCskSvyK854ja
Gb5BZfSljwFAVdS3B52IJa8qJ1ymSxOEKoDoLaxTzVOG+QAmLiC0SyAQUOUdmCZ9Z85WYAnuKwod
lMSwLABNFGPJepQMKSmkDent8VRryHTkBIBKm9hvO3gdGYyTDoUa10HtXIv0is2W28C/P+48iQiT
LXtXp9nbJ1XutUD0P6IClgtGzeEBXM09u55ltAOcJZGSnJZkA+1zApNmxzbd0NlL6tOMufrKsSf6
V3QcizGfATuBpxq0QahlkwE3XEBzlKEHbn3g/nUl12iaXDNhYVg1sbWu5U0TOLYtCy4Ki2rIKLyC
GYGPFvbHwDiOaMR7cUZlvnE4kuNOfKBfGuXpCgYj5715I0q5ouS+OJlPkR3yocd1a2Dr0ZFvKshn
m6mCTwuQhQn1VZBhE/FTuortUTzzgdfO7UuuNN2hdCc3t7gZJP4YUSpwzmO9ei0Qtc/E6/WPAzmY
aGMQ/9RCAKiOsBv8Zr1YXgyKt+wtZfihfgYnrUCvd0sKXlxy9rXSaLfBQi+xmN4PuCfEjZjuJm1U
FWstj3x/ytNwzAXVe9Lnfl3INQMYA1ZreRJyJqVoTlgryxaMegZbZHJc2JrBAUlNyog9YSfhrSXV
dNjjai0WIFuB9xhDve8OW9gPGIsiH5sFkCv710sT+gGuGwwq3/OZqfDSTdG+VKgnwNtu454m9JzS
pqxIuNvT/xTArkReEfbAnng2FnXYUmf6yY2UxSIyed5S2W9Dc5CFpN/gmj5iN4caObdZKEkarD3T
ERKDG5wlqm+GJRHm/YmmBeEAQv9fyAH7w9zEamoTxf5mvW8GRSU2jJLYIiR0a+G4E/z/oDBAxnkd
Ct3p3mjCSN0vydfvvdTflWRqpIXhCN/G8F7ULAmVXx3o/iYa5kmMgo4WSLvHVTCfWh1IGotyLh1k
XduwbnxQhfTaXjSivo+UCuOAup3ihEkhC9C1o5qLqYOv8xSjRQ6KcsH34vifyqQiGjD9bhrRJk7+
Kvhqi19Qkb94ViYiI5EMBJ+BWs5ET9OXWnjaEgGP8smMJdKBlY6S/HZ55VX8hg8RiI3hJL5AilF1
DJ2AripzAr8ux4dV+vgR4r0MlHxNMplF2JO+LF9vVVP+vj1cArQyqAA3szf8/P76zzlQBk6PJbX/
ekhPWjA5ZxdvaaO2NKZB9xzcaSs9y/fjgcTphCvIZS3EeiMtORXd9pPGXFfzt9a1btcYK+C1Cnhg
tOGROO7UsQYmtPB8crk0/iQPcgzkwlEFhNl9vT85YmLjAXqG/S+0TkHDrhBkFFUgVLDyliRz+XWc
DAltv0fVeuX0Xc+/cXfqp7oPdi5yS95Zz+S6m47qiIPXaE6WOhpxC/A/05lxcNiAYyG7YE3TlH6b
9A5PxxWv6RD77GP8JKtuw5EqWM/NxGMc67qukjfINhzWblrw0rfAl/ijqybKKDVnSGEeruPTYpYl
AbYbsXqxXlWGrrZDHdgXmDh6VytUlWU/7wkNnls6pl36kryAxG+2l5FnjgiXHFJalSUz1n2QfeNj
vGmU4tumL5c3auEPdh/C6GOxgkpkuYEYSw2vJP2E+bgxXyY2kMkC8oOrNsCJ2tfBk/qvxtZ3VXas
JQy8zTbZ6+pCqTyLb2oJhoP/0hAfmUdNCIJDBl3osYMPeF+QivpJqiGSGYkr9Z01eHaC3Zf1xwjv
BptlPe73EXs334pVRwa3OOMuPj7XZhFF4DTYp2H5WWKXAXTIwPheDRq9RaW7q+0409yGQ9pUY+1e
Evw92ZKEW6oeqXaUtH6w+7pJprH3VuUHLUU/8LsJOr8biFydzTZ/r0hN/gOIFwe4rgcEMQKgy9w2
cFiOhk7G7fQz+DwXrfyxBYZ2HroWDKoA4f9hfDyGrKg1TWUK5K5Fh9u0R4DF8necsuueb/cnOmL0
tVLyoROXgZytGCE8BEeSww0SQ7D9vpzEU8AkV1pDNZRCwHR3qmzuf5D01zXBEqg+PBbzdYHuOPT+
q8Td4iXOP95nTGhL8xQGWVU41ClNZOeb+bW3wyPcIbJ4qOxN4fqpbJIo58pN3Q/h1KNZsvzP8iRO
/TmHl6DS3zCmDtwgaRzvVCXOINqamHQrSDfgc9ho3saLT+vv76Hh9iR+0083FQ1YUN6f95JG5JnL
uq071/GzuWqXGE+WJkBdBAgpa5hHkT+gDyY2gFJcsBjliuzI6YzDoGaN+FHrI2YYodpPU8wY3BZH
ndPYpTOeylW2xZmO2D8naiCIxLgxpm5qrkzN3TRFH5E6FrjTmx64V+2XTNsKt/ArAujsiJiY6rKQ
VM5qIzVEPAkzFZ0JlEprE//OhnWHdwV7IEzzhU7JhUjLAsSctQV1tWvGCKJl86VvGA2FN4PpZK8l
FJaG33BJ2ERZ4VgtA/D00blYqvtotBfxxcnha8quv1EO/mjtB+4yCWpbPtTA2IQChoPFyyWvGk3P
m+m18zlKTsOcGc0/YHsF6zcFXpVACZMUxCJn/zkVSnHgsaj6wBoew5zM3Knqwcs6q3Q7Bt+HIVtC
PPqkReCDFKl9P4EK5G5ZXzsBwaecyFXc8oI6d+b7yI9sDs7zuOgFMO6vJe5YKunxv8xszIwxIXyp
oRddA9szpUprC0PuINJwfVmRifH7siGOSyAa3McW4Vjv6l1bLPFL11XkV9MXqPFEQ9MyyK71+Ikr
eCDrx8xiuBRHUqqbmuxH/KoL0+nzWcxu/Gn+lDGbGRE0c6KAvQorUYIjpxUM1QTzz6tGYY9o5Qm0
UWC1pQ6kcKqK9olSnUm4I6o1O2HER0kjRYoB8H0ZbZbynmpduoacVcWAUyYzw3MWdAj4+TSRQCay
vKa7cCh/E31ys1nzGUNfUo2gUYXsNOFrCJ/Eup99mHsIhRxi7fOKC1fYpGNT4J/3938FgFPyQxR3
9tduqbmDIKarj12MoWu9kANLBjuzrexwMmn4aE3NTO1SMdFqKEUH+HNM4Wj6Q9Sqdase6sqkJ53A
/yAqz1mYogeJKJ5KpZFEQWyvujeALE+1faJ1VsNYctC74T3vsEx41+YeXlaFVpLIDSHUxs18WbTz
0CXR8Iu5Cfj/Us1ciMdCHu4gW35WR9xtgWNVlrGEZLh+NciRLM0n3kW+oLVKyNfzbr7JlVdPRl/H
9BCMXhtBo/BNjboPwn7Nndo3sLm2yqDHodyq2Lhc+LfAmJOiPisgAzbqJT2Htg53uSCju+PWSuLz
CcPKIxsSiNbcC35VdXYW9GxSPmMsVfoVLzR6j6b7+a1Ctshp5R8n/nyFu+pT8deFdHEKCbSub5g9
RQGxqGoyJZKIOcfMM60v98oqFZ+D2WiCrLz9b2mRDgcBRh0/QbVCYdIRmSDKbFlPyOWimqkuv+Wh
KEF9JA8lXBhOWiM/ucA4WvtYw4YOv56vhCI0+brFRjG889+cMKILu9FLqch5CEbj6vYfEPg/2nso
ooV55ihUtfzRnF/XgZ31r75ktl/orK4Pou2NAIa6Jpt7mjSlwNY0qbURLW2dm3JV+Duvl50FIlAo
bESRSigiLm/gaae/Nv+UEzEWDYSsJqSrw8OacCqVx3knE5v8ZqTus956XBmJxX8693oUTWqFeD7x
8IKcJqDRcT2etzDJYNr3njuL1ynWDQjg6mLt1yrk2SyA4aI4Rg8NkI2iDv4UeDiR/Mj+so5dW2tX
jAH9YEbbArpU0hiKLx8R91/IOyRufthMdyGCbj3dT+2Ml3suGdTVHN+I5jenEM0wikWinQqYz+lj
opoczEnEu/zK8OddTEb2SLoJKbQ5IqzC33krByRj5phP8CGz+yQBPhzWyCF9vTnyrEN0cYSH7DvS
K6ikRHJO6HC2lcn3/ZC5oxIC8/jy68+mwFjhTq0FL/n2XRNfL+Ffi2m842MZKtuemN8Bds7GrBL+
vqepxukBsMBBRxkT7ssfS59bRLDN1lyU/bxcnI0dcdnKZiOvcY6S8DXqJ+QqeWImy1DhQgyFtXrz
kW/z4GoeLsJx+SeH3KRbx6K+sFdncA86wym+WH7OMBKPxxkwT+SgRb74YDlkDHLf4OeAMfLiPY7s
8oG8RabefqUWKCW2ITsUkM26LKDF+TsLeo659fDzXJFGefa2IPn2XgaZRFCFqtHRs1q6y6g8TcTY
t7u4BT59Opr0mc4mgjCrOgchWLMCp8IKykCa548c4vrweTrant4Wc/4vSNW6lLonzGfyjP0towKd
EAU/JPdJvjoAIuYP5pbS/a210oy1NqTknZpXfsDiWO6vLkUovcxDJYC5bwxbQ4rjXO5R77x2KsmU
mWKxd3mx/ND7uw7EjKL/6KonbXKt2WTyQ32gl4BuKNdDjHaZATYHE52JkFInl24ASgmEWV0aPLhQ
huD4GhHe4iVQ8Gl5++26s42EsPcSF8sXMy420tkDhfWdD931uoCdKE4AzvNW0zJzARcRxtfbvTtb
DtIzOHpAbgyc2QbfBxh8ki6kS5d2vO2y1GE8B1CMY0burTg7icHZUUDfLJg/a2Adr4OR5VPBP4NN
2F9gF8dA9/wsiVFfBBT+6IhKNXKR5V1E0HKGWehMGnamOevUH+7znJveSEYHA0U6xvZMNCXP631z
TJ/z9dqLkEB938ezLe5mLWQdq4y2a1gAwXvU7FHtXBUD+Ws5ZRpBBAutwcnvfQb17bwCKRRdoofQ
+0U3Ng+EdPKwdYZ8tdPaJgu7m6sGV/Ma8N+2yARldSpoWnDs+R1dalRhQixczE1irnqYr3sCRWdg
lxaSFmZ0nCGZwCb6nAfQ7TaH+iqeAHcqcUjLF9xtZR7uhctBS1SG6iShf1NapiyrgOPRXNZYlBS8
auRc787IusVFH/ixWg9wkbpBh0EkPdq40CM1UHp5zOuXXHH/+q2OUkjj+WQxJg90XhsuSiElW0Dj
h5DHMECb9ItcGLutT1uh/DhNRMLMTIg1RIFg73PwFhvYR2qIy685MSlK8DLL+bs0qVT3cJbxySiM
w34rR/q92qvxsK7riljK0omxeA5NHSzH6wMcXvDFjEn1L1Vi3hrKas4hpDp1XSoaL51PlsIzV535
6RTrQ6r6y40DWFcBcU3ss6qBZlWqXrmJ8E6R6DPLy/rUKY8kGqcW3fDsbgbevFZIaL5fwpuk5RC9
IDT2+59/e7PfZPn+8Q+6de3Eoa3KlW8kBB/ZI0+Sxl5iFC0NBQtTHlxUqxbaOd+F99Z+K0U8utRg
dMK0+903t+J+rYSlKRdaJsxF0IdVepvB+2VJqR+bdSVTRLIoA4P7HAkDyk/KieiFPRMVcjw3Iqk3
ix0cPTsInh2Cj3lp/AofReyPv0pWmCLcRiwl/xz1hV7Ii9YNU6H0ZcDKfgc2iFqMPqOgO8MALfkm
ZXS2UBebTU1/DzmJyvdNvubuPGdiHQ6f4MjSUeAO87x5KD/nOEmJn0RVLaUMrVn8oGM0jLxrJDH5
05vxwaKTJwrp4dPZDgPGubRXEGMDVDoBFBJ6Df+uNt9qBNpXrp2TYHEmGG88xOsJJJAGeqM3ptqN
rN2voaEXqptYzvSfgh2903ovIA3MUo+3/Dj/FqB8IcDjcsP9ecc2ao+2QY6BwwSaWRQedotNWdRZ
TdU8nTEK/ifxbVO6YiNfDGq9zDWNGODLVMLsuXPIPQKFCMdo854MCR21tw+izOnzUvHao7ldls13
zgnh/XHDh546eJMDCfZIwEPJPxF5FoSwUrXa5KolNKZtT25Hsp5U3wRkqrd39IjAgsqY/dA/Q/Ib
K/D26pzBjPAoGgG+UjL6nJnf66t+NF4TupOc70lN7GhI8agyxiSsjSkBu7wCIXECcwTL1/bmVILt
UO0dPCrdsaDuoZ7Qo8NFKF2mDRrozNDOR6Nvs0MthA6vYXCHDX5ZpsyFeGDyBehUTQyu6infsC8R
Yy9mQ8Eq0VcDttmZCuTMOhYbzm6bNZ7csGK9ZAkDlJdih8chc58YuEZmAYvAPrBx7xIBwJnjz6Wr
kxlV+JLTHCDt1bPB+Q00DWmXedYGkZ6oQ0/Ppt5OtZCYD6xiqIncMKOI+Yn15lBKz35La6+CRhEk
dQkPGlwDumYy2w2rxUyvC6c6p6Xl9hO5/xbExTgUrRTSLM8GBt+nck09vk0o45fWh0YRDTcO0JO2
I6coMBJS43Jmo0EbTNb4IKtTG/J1opdeZAfdxmooclDMsL2v6W1MZH3+pMt/OarwnEjnKg4q4M/o
rnczavV9udp0NMjxG9p/wvwUP2FiAtUPIY5QbFVFTOSvS/muZi7ONJHqhOE4b4b0agPbULtySJGC
/0W8GZ+bBN3XoDR7xXfpt9zAbBMmcnDjexJeev0LYqaTiw8vt7jpK2rnpCs2K8gjPbxGpNPaiMHi
aAPSnL7r489Rzb/7cfe+ryHEKn2AUnrCN1CYt73UekgtNOndGqXA9xIlou9DXTTt+8sdpfqBGugK
ASN73PXQ7EMnfLd0nm1xA4+HTN8MqW2eHOX6iihEKKCaM1iqnC1V/BQfiZAK7fP0fv7UT0QvnnFh
gD5Z4OPIZ9eQIi/kyuB0nZzfMteV4HVRZjAQe1hPuQ+IQP9sPMIUPb2FTAw8uzsKKR8N/iKmRWhx
mGoV+l6UUx1KwvLLus+szNz7jneFEN6DV8MxYnbhpSm7OrXD+r6bTxFaqeAOhp77IFmi92TXfxY9
TP/IOdDm6OY90jCsGvu9KNnSRwp1cfjpES7RbVIUz5d9wYt0xB+1wSF+DcOL/fg1EnzF1vbl2gmd
ebTtQow02sDWSoaMadpDE3iwJig/qpnMbOKMWVfLqzOQekOHtK+fGkjURoSuoof5sV3k2hDsVENq
AinjhlkTFVCOsUbh4KMTPqQqPj99JOMShGW6V+0tRomHsqwK7nyhZilGyrgXNCFLJZ9Xu2Nm6ohy
mvt629WBmppUtXJ/jVIaKISaOwUey7sPXnHmqliAjjjDv3QNHj1+bIVRDd1Z9Mc6H3JFwmFcVOCy
T+k57OKt1Nwq4Bo86RNU5mxNC+Fb6/LEJy7UjVVSZqaCE1hyOFBcBBaN8yb3K00Wt/XIXbiYIJp0
KF1WYyDG72wDUY+7RqwqL7/eB/poS8KsfWQKyaCbS4NvFMmfMspq5gjBzD15hLxbpjjQsG4wo37O
HOTkEbQPr0QUFiwA+kmAoUm5yTpsplpwVzARKPgwhdZbeWY10zYM8dDy2xYfx85Rg0jMXkrqsTQV
OmQ1awQGSNHns8+3q3/arWv9eGqP8f0qxitwNwSN6zWzeObbTsIS0qO6D60FSOTHCWtqjfW7tGAE
MOb5qvDjSPdcj35/Ai+ezE2Jv+dCn1ld2inKodIVVZB22YPp6t7Hm3RObbtISjqGEkDeSfsMjzMd
hLYK6fr+OWwGF/wABcs6PjZAhSTEbXZekY98m+GogGPeHrdeRFRf3JRCThKpUlj1GiknwQg4D9e1
YghpxOBCdudTHL95P97M327QCI1UFi33h1NUuBxnWl2u4k92US8spPrUETBI2WpYaHd2NZuZQabv
HtIizD/3/a+L9MIg5dI7n7HqSqfQNWBlqzcz37RX22678JQlYpj/j804Yopdc3hEHQ4UxDAPFrEz
rw90n2Y2lSonoKN8fBCgxVJP7xogsNrLYEgw2oAOIGVkyAT6ZmLsu0WFZh9u0+aamLQEcmgaS9G0
JQEZZPxscKrB7A9eeeXhYwxs/ExK5g9PyC32kgE+qdbNWfo4uqjp1bSBLvLn1xPFPZE/bavpFk40
uCbcLVWn2YQ7nFwsOTPM3jYOPVwcjl/sv9nFbTW86XqY9Y3TiMzDJyGe6tjUxGmUo6T7YFkIIfsc
WyAD1zmNOYtbOBdTXWg9/QhVyoH1Uz9m+flZmiMfDxUqxJD1hihLBWshHeOCHSAzTVN7XYhlPIUQ
MZzGpTKfEZS1aB/T55fS9Twn+y1JcO/xQMNCg33IjCQofTyQlnyM9G/8IosQNioX2qYb5fD3vWiY
TQTPcgVAXqXlLkwOPAZ9y4BQ6OnvSN5wYjIgAFPxx9WXDM5AlRgMsZ6zkQ0G5Uw4oPwACLC8T2p1
srtIi8BLiITSQ8JyM7l7+DzZ84OlSKRpaOb4h6hnkZiTyCeGwVNwazoJ+VkTYS9PCJvaQw6XsaXD
EJ8aYunuJNlHw4bWdwjXRpgdHT+UK+i5sqoUtToyNowT1ApszPvWgyjGMk8cZelV2kB658znP96g
u6zXfXOhOwgpY7rwoYAqbYfW2VWWL2oZb09l+bBhOI9v2pbXm/qiJ/bGybAiT9eIlbJaUrL/klTm
8j2uZg5Ur5vGxfZe6pC6WEhQxkI7Pw3p6uEOpZw9Bi8A0pIuRSytqH4u+1ufT2mTmcMSxxWjABMg
ELlV+IUgqUAYH1bb+lF8w/+KvA109fJPhcHLSF1SN5xhvlYwn+cdTtxdTd4gdT/WijR0rhWTnYik
Z/7q481JRA2bJe+F659X+F9404N4nkkdSYkMS+Rwwqik1ReqQx2wa0wEoK+tWqFZw/fQJTDjEhaw
8j7QNEx3RojRdL8V2Zu+j506nBN/6hShGlQy3T8YMEwTPrx4zi9wm0CRU99Wjmw1XIdQ4b74ucZR
/egQT5zRhZZHQEirOG/Az2JI2PVwPxqj7+84HspIwhxvPEVV4m0Y1LLin0XEIQ26GZiRfVChHU2t
O/xnd7hsRcWzb9HafMPVorlwywRUXB0DtM1mVowctXPtNeYkxTdyiSuh9ssHpWsFoue7PW5hGoyi
0L//8LQqM9cbgl/HSqcPCKh/M6oet4FrXo1Nc83/C++Kgyxth5jxA4dLQPGvB7rdLZCq81mIuhAg
EnJt3F69MGTuyxgA3D6RKOW/cf8S5Ri6sWtEjJ4C5FoYPGGI4jv/FoIOLJ4JQxRiKiV6F+8h1snQ
BIzzZmQHr0L4P7Ix/CimW+CeZ1dXkuKuZoGr31Prm3zpLQhwMwwWeGAcFpyHyVDsr+5VW8cIpZ2W
2LoLCP2/gnWY2gDNBSUwkAmhtFUznap9KuU5pjmMb2ZqARdi/HX19gvqfl/1YzOZe54rhZ35+dyu
dwWpcsXM9rHJ/U1s4tnGns0Z0fmED79P2mx8g1QrKbmbmcjhD1rCvCMWARWKp5lcRm1Qq9f+BVOW
j9xlVbs1lx6I7omtO9fGL4mdy34kpOmrTUETDI9pReZb7Z5gnawIGrTtYQJQ5DtM09tyFn/5Wf5W
qIx8gzEv4qMFmQ7hj17YMvn3wJuUG1M2muNYhiOsx79QLU1OXatDFPYkfDi1vY5jURb3+/hn5Sqd
cd0ncy/tHXBKgMS24hfLSx9yD6cecz1RSlB5ikt1PUXmhoXGJHQCSOOUK9K5+egBRRuDx0nKwMLC
TZJ09gkRWxQh/lKqsw3+IWYCh1od7Xc8MzA/0resNNqa8935bRz1kzsBoUBC4TxVx7fJrmGCopG6
GYLQF2u5cJmQeN7WFo0jGz4y5uwMOh7W8eXhyhGyBvM99/H+WLDKtMxyoSXg2IAExceIzP+peJKq
ZSEBnsfWd3SZQvKM91iQAzBURlQ2Bxg4GsoqSsi3d8wFAajQ7RCjXe06dckawrf7Yd4jF+DYpldu
ZgJRD32ZcTPnTeydFPqEbgyEQ5pI//kRVKtYV6LbJnWtgDbSY7QQ7UbD2lIsMNaZ084GX8l4HClC
H6ki9tYd2v5BN47fJDXDnzuJ1ygud8ldoX3zWP1UARvs62g9b3V54AaYwlVUFNGebHLQRwBxDAEE
+XESBmPyNHiAqNnZYQNGccQFR+sK7fnSl9m5Ah2igBfeFDKB+qKjIicDwy+fCBVbpziM1RBbevS5
j+9Kb5FDVOo17dmzoPAitUG4tAu7JD07+z7xNHTZ2i+Q+Fo5HRDOpQVFt6tLrVAVpJraWujW1CEn
5dV7gGX3R/rweoBUBec4k6NYmpN9fPRN9o3uTcGSbDTRsRALH6AU3bF7kqLgeAGbbTYM+0oDs9kp
qFX3QLSS
`pragma protect end_protected

